library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ControlMemory256x42 is
  port ( In_car : in STD_LOGIC_VECTOR(16 downto 0);
         FL : out std_logic; -- 0
         RZ : out std_logic; -- 1
         RN : out std_logic; -- 2
         RC : out std_logic; -- 3
         RV : out std_logic; -- 4
         MW : out std_logic; -- 5
         MM : out std_logic; -- 6
         RW : out std_logic; -- 7
         MD : out std_logic; -- 8
         FS : out std_logic_vector(4 downto 0); -- 9 to 13
         MB : out std_logic; -- 14
         TB : out std_logic; -- 15
         TA : out std_logic; -- 16
         TD : out std_logic; -- 17
         PL : out std_logic; -- 18
         PI : out std_logic; -- 19
         IL : out std_logic; -- 20
         MC : out std_logic; -- 21
         MS : out std_logic_vector(2 downto 0); -- 22 to 24
         NA : out std_logic_vector(16 downto 0) -- 25 to 41
  );
end ControlMemory256x42;
-- FS: FU_s ALU_s S  Cin
-- FS: 0    0    00 0
architecture Behavioral of ControlMemory256x42 is
  type mem_array is array(0 to 255) of STD_LOGIC_VECTOR(41 downto 0);
    -- initialise the control memory
    signal ControlMemory256x42 : mem_array := (
      -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
      -- | Next Address | MS | M| I| P| P| T| T| T| M| FS |M|R|M|M|R|R|R|R|F|
      -- | Next Address | MS | C| L| I| L| D| A| B| B| FS |D|W|M|W|V|C|N|Z|L|
      -- "00000000000000000 000 0 0 0 0 0 0 0 0 00000 0 0 0 0 0 0 0 0 0"
      -- "00000000011000000 001 0 0 0 1 0 0 0 0 00000 0 0 0 0 0 0 0 0 0" B
      -- "00000000011000000 001 0 0 0 0 0 0 0 1 00010 0 1 0 0 0 0 0 0 0"
      -- "00000000000000011 001 0 0 0 0 0 0 0 0 00001 0 1 0 0 0 0 0 0 0"
      "000000000110000000010000000100010010000000", --0 ADI
      "000000000110000000010000000000001010000000", --1 INC
      "000000000110000000010000000001100010000000", --2 XOR
      "000000000110000000010000000000000110000000", --3 LDR
      "000000000110000001110100100010010010000000", --4 Sr nB
      "000000000110000000010000000000000000100000", --5 STR
      "000000000110000001110100100010100010000000", --6 Sl
      "000000000110000000010000000001110010000000", --7 NOT
      "000000000110000000010000000000010010000000", --8 ADD
      "000000000100001100010000000000000110000000", --9 LRI
      "000000000000010100000000000000000000000000", --10
      "000000000001010101000001111010000010000000", --11 BEQ
      "000000000110000000010000000000000000000000", --12 Catch
      "000000000001010101110000000000000000000000", --13 BNZ
      "000000000110000000010000000000000000000000", --14 Catch
      "000000000110000000010000100000101010000000", --15 CMP
      "000000000000100000000000000000000000000000", --16
      "000000000000100010000000000000000000000000", --17
      "000000000000100100000000000000000000000000", --18
      "000000000000100110000000000000000000000000", --19
      "000000000000101000000000000000000000000000", --20
      "000000000000101010000000000000000000000000", --21
      "000000000000101100000000000000000000000000", --22
      "000000000000101110000000000000000000000000", --23
      "000000000000110000000000000000000000000000", --24
      "000000000000110010000000000000000000000000", --25
      "000000000000110100000000000000000000000000", --26
      "000000000000110110000000000000000000000000", --27
      "000000000000111000000000000000000000000000", --28
      "000000000000111010000000000000000000000000", --29
      "000000000000111100000000000000000000000000", --30
      "000000000000111110000000000000000000000000", --31
      "000000000001000000000000000000000000000000", --32
      "000000000001000010000000000000000000000000", --33
      "000000000001000100000000000000000000000000", --34
      "000000000001000110000000000000000000000000", --35
      "000000000001001000000000000000000000000000", --36
      "000000000001001010000000000000000000000000", --37
      "000000000001001100000000000000000000000000", --38
      "000000000001001110000000000000000000000000", --39
      "000000000001010000000000000000000000000000", --40
      "000000000110000000010000000000000110000000", --41 LR
      "000000000110000000010001000000000000000000", --42 B
      "000000000001010110000000000000000000000000", --43
      "000000000001011000000000000000000000000000", --44
      "000000000001011010000000000000000000000000", --45
      "000000000001011100000000000000000000000000", --46
      "000000000001011110000000000000000000000000", --47
      "000000000001100000000000000000000000000000", --48
      "000000000001100010000000000000000000000000", --49
      "000000000001100100000000000000000000000000", --50
      "000000000001100110000000000000000000000000", --51
      "000000000001101000000000000000000000000000", --52
      "000000000001101010000000000000000000000000", --53
      "000000000001101100000000000000000000000000", --54
      "000000000001101110000000000000000000000000", --55
      "000000000001110000000000000000000000000000", --56
      "000000000001110010000000000000000000000000", --57
      "000000000001110100000000000000000000000000", --58
      "000000000001110110000000000000000000000000", --59
      "000000000001111000000000000000000000000000", --60
      "000000000001111010000000000000000000000000", --61
      "000000000001111100000000000000000000000000", --62
      "000000000001111110000000000000000000000000", --63
      "000000000010000000000000000000000000000000", --64
      "000000000010000010000000000000000000000000", --65
      "000000000010000100000000000000000000000000", --66
      "000000000010000110000000000000000000000000", --67
      "000000000010001000000000000000000000000000", --68
      "000000000010001010000000000000000000000000", --69
      "000000000010001100000000000000000000000000", --70
      "000000000010001110000000000000000000000000", --71
      "000000000010010000000000000000000000000000", --72
      "000000000010010010000000000000000000000000", --73
      "000000000010010100000000000000000000000000", --74
      "000000000010010110000000000000000000000000", --75
      "000000000010011000000000000000000000000000", --76
      "000000000010011010000000000000000000000000", --77
      "000000000010011100000000000000000000000000", --78
      "000000000010011110000000000000000000000000", --79
      "000000000010100000000000000000000000000000", --80
      "000000000010100010000000000000000000000000", --81
      "000000000010100100000000000000000000000000", --82
      "000000000010100110000000000000000000000000", --83
      "000000000010101000000000000000000000000000", --84
      "000000000010101010000000000000000000000000", --85
      "000000000010101100000000000000000000000000", --86
      "000000000010101110000000000000000000000000", --87
      "000000000010110000000000000000000000000000", --88
      "000000000010110010000000000000000000000000", --89
      "000000000010110100000000000000000000000000", --90
      "000000000010110110000000000000000000000000", --91
      "000000000010111000000000000000000000000000", --92
      "000000000010111010000000000000000000000000", --93
      "000000000010111100000000000000000000000000", --94
      "000000000010111110000000000000000000000000", --95
      "000000000011000000000000000000000000000000", --96
      "000000000011000010000000000000000000000000", --97
      "000000000011000100000000000000000000000000", --98
      "000000000011000110000000000000000000000000", --99
      "000000000011001000000000000000000000000000", --100
      "000000000011001010000000000000000000000000", --101
      "000000000011001100000000000000000000000000", --102
      "000000000011001110000000000000000000000000", --103
      "000000000011010000000000000000000000000000", --104
      "000000000011010010000000000000000000000000", --105
      "000000000011010100000000000000000000000000", --106
      "000000000011010110000000000000000000000000", --107
      "000000000011011000000000000000000000000000", --108
      "000000000011011010000000000000000000000000", --109
      "000000000011011100000000000000000000000000", --110
      "000000000011011110000000000000000000000000", --111
      "000000000011100000000000000000000000000000", --112
      "000000000011100010000000000000000000000000", --113
      "000000000011100100000000000000000000000000", --114
      "000000000011100110000000000000000000000000", --115
      "000000000011101000000000000000000000000000", --116
      "000000000011101010000000000000000000000000", --117
      "000000000011101100000000000000000000000000", --118
      "000000000011101110000000000000000000000000", --119
      "000000000011110000000000000000000000000000", --120
      "000000000011110010000000000000000000000000", --121
      "000000000011110100000000000000000000000000", --122
      "000000000011110110000000000000000000000000", --123
      "000000000011111000000000000000000000000000", --124
      "000000000011111010000000000000000000000000", --125
      "000000000011111100000000000000000000000000", --126
      "000000000011111110000000000000000000000000", --127
      "000000000100000000000000000000000000000000", --128
      "000000000100000010000000000000000000000000", --129
      "000000000100000100000000000000000000000000", --130
      "000000000100000110000000000000000000000000", --131
      "000000000100001000000000000000000000000000", --132
      "000000000100001010000000000000000000000000", --133
      "000000000110000000010000010000000110000000", --134 LRI2
      "000000000110000000010000000000000000000000", --135 Catch
      "000000000100010000000000000000000000000000", --136
      "000000000100010010000000000000000000000000", --137
      "000000000100010100000000000000000000000000", --138
      "000000000100010110000000000000000000000000", --139
      "000000000100011000000000000000000000000000", --140
      "000000000100011010000000000000000000000000", --141
      "000000000100011100000000000000000000000000", --142
      "000000000100011110000000000000000000000000", --143
      "000000000100100000000000000000000000000000", --144
      "000000000100100010000000000000000000000000", --145
      "000000000100100100000000000000000000000000", --146
      "000000000100100110000000000000000000000000", --147
      "000000000100101000000000000000000000000000", --148
      "000000000100101010000000000000000000000000", --149
      "000000000100101100000000000000000000000000", --150
      "000000000100101110000000000000000000000000", --151
      "000000000100110000000000000000000000000000", --152
      "000000000100110010000000000000000000000000", --153
      "000000000100110100000000000000000000000000", --154
      "000000000100110110000000000000000000000000", --155
      "000000000100111000000000000000000000000000", --156
      "000000000100111010000000000000000000000000", --157
      "000000000100111100000000000000000000000000", --158
      "000000000100111110000000000000000000000000", --159
      "000000000101000000000000000000000000000000", --160
      "000000000101000010000000000000000000000000", --161
      "000000000101000100000000000000000000000000", --162
      "000000000101000110000000000000000000000000", --163
      "000000000101001000000000000000000000000000", --164
      "000000000101001010000000000000000000000000", --165
      "000000000101001100000000000000000000000000", --166
      "000000000101001110000000000000000000000000", --167
      "000000000101010000000000000000000000000000", --168
      "000000000101010010000000000000000000000000", --169
      "000000000101010100000000000000000000000000", --170
      "000000000101010110000000000000000000000000", --171
      "000000000101011000000000000000000000000000", --172
      "000000000101011010000000000000000000000000", --173
      "000000000101011100000000000000000000000000", --174
      "000000000101011110000000000000000000000000", --175
      "000000000101100000000000000000000000000000", --176
      "000000000101100010000000000000000000000000", --177
      "000000000101100100000000000000000000000000", --178
      "000000000101100110000000000000000000000000", --179
      "000000000101101000000000000000000000000000", --180
      "000000000101101010000000000000000000000000", --181
      "000000000101101100000000000000000000000000", --182
      "000000000101101110000000000000000000000000", --183
      "000000000101110000000000000000000000000000", --184
      "000000000101110010000000000000000000000000", --185
      "000000000101110100000000000000000000000000", --186
      "000000000101110110000000000000000000000000", --187
      "000000000101111000000000000000000000000000", --188
      "000000000101111010000000000000000000000000", --189
      "000000000101111100000000000000000000000000", --190
      "000000000101111110000000000000000000000000", --191
      "000000000110000010000110000000000001000000", --192 IF
      "000000000000000000011000000000000000000000", --193 EXO
      "000000000110000100000000000000000000000000", --194
      "000000000110000110000000000000000000000000", --195
      "000000000110001000000000000000000000000000", --196
      "000000000110001010000000000000000000000000", --197
      "000000000110001100000000000000000000000000", --198
      "000000000110001110000000000000000000000000", --199
      "000000000110010000000000000000000000000000", --200
      "000000000110010010000000000000000000000000", --201
      "000000000110010100000000000000000000000000", --202
      "000000000110010110000000000000000000000000", --203
      "000000000110011000000000000000000000000000", --204
      "000000000110011010000000000000000000000000", --205
      "000000000110011100000000000000000000000000", --206
      "000000000110011110000000000000000000000000", --207
      "000000000110100000000000000000000000000000", --208
      "000000000110100010000000000000000000000000", --209
      "000000000110100100000000000000000000000000", --210
      "000000000110100110000000000000000000000000", --211
      "000000000110101000000000000000000000000000", --212
      "000000000110101010000000000000000000000000", --213
      "000000000110101100000000000000000000000000", --214
      "000000000110101110000000000000000000000000", --215
      "000000000110110000000000000000000000000000", --216
      "000000000110110010000000000000000000000000", --217
      "000000000110110100000000000000000000000000", --218
      "000000000110110110000000000000000000000000", --219
      "000000000110111000000000000000000000000000", --220
      "000000000110111010000000000000000000000000", --221
      "000000000110111100000000000000000000000000", --222
      "000000000110111110000000000000000000000000", --223
      "000000000111000000000000000000000000000000", --224
      "000000000111000010000000000000000000000000", --225
      "000000000111000100000000000000000000000000", --226
      "000000000111000110000000000000000000000000", --227
      "000000000111001000000000000000000000000000", --228
      "000000000111001010000000000000000000000000", --229
      "000000000111001100000000000000000000000000", --230
      "000000000111001110000000000000000000000000", --231
      "000000000111010000000000000000000000000000", --232
      "000000000111010010000000000000000000000000", --233
      "000000000111010100000000000000000000000000", --234
      "000000000111010110000000000000000000000000", --235
      "000000000111011000000000000000000000000000", --236
      "000000000111011010000000000000000000000000", --237
      "000000000111011100000000000000000000000000", --238
      "000000000111011110000000000000000000000000", --239
      "000000000111100000000000000000000000000000", --240
      "000000000111100010000000000000000000000000", --241
      "000000000111100100000000000000000000000000", --242
      "000000000111100110000000000000000000000000", --243
      "000000000111101000000000000000000000000000", --244
      "000000000111101010000000000000000000000000", --245
      "000000000111101100000000000000000000000000", --246
      "000000000111101110000000000000000000000000", --247
      "000000000111110000000000000000000000000000", --248
      "000000000111110010000000000000000000000000", --249
      "000000000111110100000000000000000000000000", --250
      "000000000111110110000000000000000000000000", --251
      "000000000111111000000000000000000000000000", --252
      "000000000111111010000000000000000000000000", --253
      "000000000111111100000000000000000000000000", --254
      "000000000111111110000000000000000000000000"  --255
    );

  signal adr_content : STD_LOGIC_VECTOR(41 downto 0);

  begin
    adr_content <= ControlMemory256x42(to_integer(unsigned(In_car(8 downto 0))));

    FL <= adr_content(0); -- 0
    RZ <= adr_content(1); -- 1
    RN <= adr_content(2); -- 2
    RC <= adr_content(3); -- 3
    RV <= adr_content(4); -- 4
    MW <= adr_content(5); -- 5
    MM <= adr_content(6); -- 6
    RW <= adr_content(7); -- 7
    MD <= adr_content(8); -- 8
    FS <= adr_content(13 downto 9); -- 9 to 13
    MB <= adr_content(14); -- 14
    TB <= adr_content(15); -- 15
    TA <= adr_content(16); -- 16
    TD <= adr_content(17); -- 17
    PL <= adr_content(18); -- 18
    PI <= adr_content(19); -- 19
    IL <= adr_content(20); -- 20
    MC <= adr_content(21); -- 21
    MS <= adr_content(24 downto 22); -- 22 to 24
    NA <= adr_content(41 downto 25); -- 25 to 41
end Behavioral;
